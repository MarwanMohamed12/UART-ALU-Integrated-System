module Rx_edge_bit_counter ();





endmodule