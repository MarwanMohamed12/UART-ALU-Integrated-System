module ANDX (C,A,B);

input A,B ;
output C;

assign C = A & B ;


endmodule

